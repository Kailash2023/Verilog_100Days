module Bin_Ex3(
    input [3:0]bin_in,
    output [3:0]ex3_out
    );
    
    assign ex3_out = bin_in + 4'b0011 ;
    
    
endmodule
